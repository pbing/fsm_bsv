/* fsm1_pkgs for abstract encoded enums */

package fsm1_pkg;
   typedef enum {IDLE,
                 READ,
                 DLY,
                 DONE,
                 XXX } state_e;
endpackage
